# KERNEL: ASDB file was created in location /home/runner/dataset.asdb
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=1 DATA_IN=58 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=142 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=1 DATA_IN=209 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=46 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=198 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=1 DATA_IN=239 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=179 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=1 DATA_IN=67 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=52 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=143 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=1 DATA_IN=96 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=18 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=1 DATA_IN=225 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=148 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----GENERATOR CLASS-----
# KERNEL: [0]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=29 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [5]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=1 DATA_IN=58 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [5]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=1 DATA_IN=58 | DATA_OUT=0 FULL=0 |  EMPTY=1
# KERNEL: Error: scoreboard.sv (31): [SCB] Attempted READ when EMPTY!
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [15]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=142 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [15]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=142 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: [SCB] WRITE: 8e
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [25]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=1 DATA_IN=209 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [25]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=1 DATA_IN=209 | DATA_OUT=142 FULL=0 |  EMPTY=0
# KERNEL: [SCB] WRITE: d1
# KERNEL: [SCB] READ: 8e
# KERNEL: [SCB] PASS: READ=8e EXP=8e
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [35]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=46 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [35]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=46 | DATA_OUT=142 FULL=0 |  EMPTY=0
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [45]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=198 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [45]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=198 | DATA_OUT=142 FULL=0 |  EMPTY=0
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [55]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=1 DATA_IN=239 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [55]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=1 DATA_IN=239 | DATA_OUT=209 FULL=0 |  EMPTY=0
# KERNEL: [SCB] WRITE: ef
# KERNEL: [SCB] READ: d1
# KERNEL: [SCB] PASS: READ=d1 EXP=d1
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [65]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=179 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [65]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=179 | DATA_OUT=209 FULL=0 |  EMPTY=0
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [75]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=1 DATA_IN=67 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [75]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=1 DATA_IN=67 | DATA_OUT=239 FULL=0 |  EMPTY=0
# KERNEL: [SCB] WRITE: 43
# KERNEL: [SCB] READ: ef
# KERNEL: [SCB] PASS: READ=ef EXP=ef
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [85]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=52 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [85]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=52 | DATA_OUT=239 FULL=0 |  EMPTY=0
# KERNEL: [SCB] WRITE: 34
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [95]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=143 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [95]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=143 | DATA_OUT=239 FULL=0 |  EMPTY=0
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [105]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=1 DATA_IN=96 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [105]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=1 DATA_IN=96 | DATA_OUT=67 FULL=0 |  EMPTY=0
# KERNEL: [SCB] READ: 43
# KERNEL: [SCB] PASS: READ=43 EXP=43
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [115]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=18 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [115]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=18 | DATA_OUT=67 FULL=0 |  EMPTY=0
# KERNEL: [SCB] WRITE: 12
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [125]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=1 DATA_IN=225 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [125]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=1 DATA_IN=225 | DATA_OUT=52 FULL=0 |  EMPTY=0
# KERNEL: [SCB] READ: 34
# KERNEL: [SCB] PASS: READ=34 EXP=34
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [135]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=148 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [135]  | RST=1 | CS=1 | WR_ENB=1 | RD_ENB=0 DATA_IN=148 | DATA_OUT=52 FULL=0 |  EMPTY=0
# KERNEL: [SCB] WRITE: 94
# KERNEL: -----DRIVER CLASS-----
# KERNEL: [145]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=29 | DATA_OUT=0 FULL=0 |  EMPTY=0
# KERNEL: -----MONITOR CLASS-----
# KERNEL: [145]  | RST=1 | CS=1 | WR_ENB=0 | RD_ENB=0 DATA_IN=29 | DATA_OUT=52 FULL=0 |  EMPTY=0
# RUNTIME: Info: RUNTIME_0068 $finish called.
# KERNEL: Time: 157 ns,  Iteration: 0,  Instance: /testbench/t,  Process: @INITIAL#6_0@.
# KERNEL: stopped at time: 157 ns
# VSIM: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.
Done
