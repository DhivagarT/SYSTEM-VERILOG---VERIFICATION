KERNEL: Time=0 A=0 B=1 C=0 Sum=0 Carry=0 
# KERNEL: Generator Class
# KERNEL: Time=0 A=1 B=0 C=0 Sum=0 Carry=0 
# KERNEL: Generator Class
# KERNEL: Time=0 A=1 B=1 C=1 Sum=0 Carry=0 
# KERNEL: Driver Class
# KERNEL: Time=2 A=0 B=1 C=0 Sum=0 Carry=0 
# KERNEL: Monitor Class
# KERNEL: Time=2 A=0 B=1 C=0 Sum=1 Carry=0 
# KERNEL: Scoreboard Class
# KERNEL: Time=2 A=0 B=1 C=0 Sum=1 Carry=0 
# KERNEL: ----PASS----
# KERNEL: Driver Class
# KERNEL: Time=4 A=1 B=0 C=0 Sum=0 Carry=0 
# KERNEL: Monitor Class
# KERNEL: Time=4 A=1 B=0 C=0 Sum=1 Carry=0 
# KERNEL: Scoreboard Class
# KERNEL: Time=4 A=1 B=0 C=0 Sum=1 Carry=0 
# KERNEL: ----PASS----
# KERNEL: Driver Class
# KERNEL: Time=6 A=1 B=1 C=1 Sum=0 Carry=0 
# KERNEL: Monitor Class
# KERNEL: Time=6 A=1 B=1 C=1 Sum=1 Carry=1 
# KERNEL: Scoreboard Class
# KERNEL: Time=6 A=1 B=1 C=1 Sum=1 Carry=1 
# KERNEL: ----PASS----
# RUNTIME: Info: RUNTIME_0068 $finish called.
