interface intf;
  logic clk;
  logic rst;
  logic enb;
  logic [2:0]count;
    
endinterface
