# KERNEL: ----Generator Class---
# KERNEL: Time=0  Rst=0 D=1 Q=0
# KERNEL: ----Generator Class----
# KERNEL: Time=0  Rst=1 D=0 Q=0
# KERNEL: ----Generator Class----
# KERNEL: Time=0  Rst=1 D=1 Q=0
# KERNEL: ----Driver Class----
# KERNEL: Time=2  Rst=0 D=1 Q=0
# KERNEL: ----Monitor Class----
# KERNEL: Time=3  Rst=0 D=1 Q=0
# KERNEL: ---PASS---
# KERNEL: ----Scoreboard Class----
# KERNEL: Time=3  Rst=0 D=1 Q=0
# KERNEL: ----Driver Class----
# KERNEL: Time=6  Rst=1 D=0 Q=0
# KERNEL: ----Monitor Class----
# KERNEL: Time=7  Rst=1 D=0 Q=0
# KERNEL: ---PASS---
# KERNEL: ----Scoreboard Class----
# KERNEL: Time=7  Rst=1 D=0 Q=0
# KERNEL: ----Driver Class----
# KERNEL: Time=10  Rst=1 D=1 Q=0
# KERNEL: ----Monitor Class----
# KERNEL: Time=11  Rst=1 D=1 Q=0
# KERNEL: ---PASS---
# KERNEL: ----Scoreboard Class----
# KERNEL: Time=11  Rst=1 D=1 Q=0
# RUNTIME: Info: RUNTIME_0068 $finish called.
