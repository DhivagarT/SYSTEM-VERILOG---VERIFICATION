class generator;
  transaction trans;
  mailbox m1;
  
  function new(mailbox m1);
    this.m1=m1;
  endfunction
  
  task main();
    repeat(3)begin
      trans=new();
      trans.randomize();
      m1.put(trans);
      trans.display("Generator Class");
    end
  endtask
endclass
